module main;
endmodule // main
