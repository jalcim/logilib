module and4(bus, s);
endmodule; // and4

module and8(bus, s);
endmodule; // and8
