module gate_not (e1, s);
   input e1;
   output s;

   not not0(s, e1);
endmodule // not
